`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/26/2025 01:56:54 PM
// Design Name: 
// Module Name: tb_mux8X1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_mux8X1(

    );
    // Inputs
    reg [7:0] I;
    reg [2:0] s;
    
    // Output
    wire out;

    // Instantiate the 8x1 Multiplexer
    mux8x1 DUT (
        .I(I), 
        .s(s), 
        .out(out)
    );

    // Test sequence
    initial begin
        I = 8'b00000001; s = 3'b000; #10;
        I = 8'b00000010; s = 3'b001; #10;
        I = 8'b00000100; s = 3'b010; #10;
        I = 8'b00001000; s = 3'b011; #10;
        I = 8'b00010000; s = 3'b100; #10;
        I = 8'b00100000; s = 3'b101; #10;
        I = 8'b01000000; s = 3'b110; #10;
        I = 8'b10000000; s = 3'b111; #10;    
    
    
    
    
    
    
    
    
    
    
    
//        I = 8'b00000001; s = 3'b000; #10;
//        I = 8'b00000010; s = 3'b000; #10;
//        I = 8'b00000100; s = 3'b000; #10;
//        I = 8'b00001000; s = 3'b000; #10;
//        I = 8'b00010000; s = 3'b000; #10;
//        I = 8'b00100000; s = 3'b000; #10;
//        I = 8'b01000000; s = 3'b000; #10;
//        I = 8'b10000000; s = 3'b000; #10;

//        I = 8'b00000001; s = 3'b001; #10;
//        I = 8'b00000010; s = 3'b001; #10;
//        I = 8'b00000100; s = 3'b001; #10;
//        I = 8'b00001000; s = 3'b001; #10;
//        I = 8'b00010000; s = 3'b001; #10;
//        I = 8'b00100000; s = 3'b001; #10;
//        I = 8'b01000000; s = 3'b001; #10;
//        I = 8'b10000000; s = 3'b001; #10;


//        I = 8'b00000001; s = 3'b010; #10;
//        I = 8'b00000010; s = 3'b010; #10;
//        I = 8'b00000100; s = 3'b010; #10;
//        I = 8'b00001000; s = 3'b010; #10;
//        I = 8'b00010000; s = 3'b010; #10;
//        I = 8'b00100000; s = 3'b010; #10;
//        I = 8'b01000000; s = 3'b010; #10;
//        I = 8'b10000000; s = 3'b010; #10;


//        I = 8'b00000001; s = 3'b011; #10;
//        I = 8'b00000010; s = 3'b011; #10;
//        I = 8'b00000100; s = 3'b011; #10;
//        I = 8'b00001000; s = 3'b011; #10;
//        I = 8'b00010000; s = 3'b011; #10;
//        I = 8'b00100000; s = 3'b011; #10;
//        I = 8'b01000000; s = 3'b011; #10;
//        I = 8'b10000000; s = 3'b011; #10;


//        I = 8'b00000001; s = 3'b100; #10;
//        I = 8'b00000010; s = 3'b100; #10;
//        I = 8'b00000100; s = 3'b100; #10;
//        I = 8'b00001000; s = 3'b100; #10;
//        I = 8'b00010000; s = 3'b100; #10;
//        I = 8'b00100000; s = 3'b100; #10;
//        I = 8'b01000000; s = 3'b100; #10;
//        I = 8'b10000000; s = 3'b100; #10;


//        I = 8'b00000001; s = 3'b101; #10;
//        I = 8'b00000010; s = 3'b101; #10;
//        I = 8'b00000100; s = 3'b101; #10;
//        I = 8'b00001000; s = 3'b101; #10;
//        I = 8'b00010000; s = 3'b101; #10;
//        I = 8'b00100000; s = 3'b101; #10;
//        I = 8'b01000000; s = 3'b101; #10;
//        I = 8'b10000000; s = 3'b101; #10;


//        I = 8'b00000001; s = 3'b110; #10;
//        I = 8'b00000010; s = 3'b110; #10;
//        I = 8'b00000100; s = 3'b110; #10;
//        I = 8'b00001000; s = 3'b110; #10;
//        I = 8'b00010000; s = 3'b110; #10;
//        I = 8'b00100000; s = 3'b110; #10;
//        I = 8'b01000000; s = 3'b110; #10;
//        I = 8'b10000000; s = 3'b110; #10;


//        I = 8'b00000001; s = 3'b111; #10;
//        I = 8'b00000010; s = 3'b111; #10;
//        I = 8'b00000100; s = 3'b111; #10;
//        I = 8'b00001000; s = 3'b111; #10;
//        I = 8'b00010000; s = 3'b111; #10;
//        I = 8'b00100000; s = 3'b111; #10;
//        I = 8'b01000000; s = 3'b111; #10;
//        I = 8'b10000000; s = 3'b111; #10;
        
        $finish;
    end
    
    // Monitor changes
    initial begin
        $monitor("Time = %0t | I = %b | s = %b | out = %b", $time, I, s, out);
    end
endmodule
//module tb_mux8X1();
//    // Inputs
//    reg [7:0] I;
//    reg [2:0] s;
    
//    // Output
//    wire out;

//    // Instantiate the 8x1 Multiplexer
//    mux8x1 DUT (
//        .I(I), 
//        .s(s), 
//        .out(out)
//    );

//    // Test sequence
//    initial begin
//        I = 8'b10101010; // Assigning a pattern to I
        
//        // Iterate over all select values
//        s = 3'b000; #10;
//        s = 3'b001; #10;
//        s = 3'b010; #10;
//        s = 3'b011; #10;
//        s = 3'b100; #10;
//        s = 3'b101; #10;
//        s = 3'b110; #10;
//        s = 3'b111; #10;

//        #10;
//        $finish;
//    end
    
//    // Monitor changes
//    initial begin
//        $monitor("Time = %0t | I = %b | s = %b | out = %b", $time, I, s, out);
//    end
//endmodule
